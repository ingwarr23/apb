package apb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_config.svh"
  `include "apb_seq_item.svh"
  `include "apb_driver.svh"
  `include "apb_sequencer.svh"
  `include "apb_monitor.svh"
  `include "apb_agent.svh"

  `include "apb_seqlib/apb_read_seq.svh"

endpackage: apb_pkg