package test_list_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import apb_pkg::*;
  import top_env_pkg::*;
  import seqlib_pkg::*;
//  import adder_4_bit_env_pkg::*;
//  import adder_4_bit_seq_list::*;
  
  `include "normal_test.svh"

endpackage 