package top_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import apb_pkg::*;

  `include "top_env_config.svh"
  `include "top_env.svh"

endpackage: top_env_pkg