package seqlib_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import apb_pkg::*;

  `include "base_seq.svh"

endpackage: seqlib_pkg