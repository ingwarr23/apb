package globals_pkg;
  parameter T_APB_CLK_NS = 20;
endpackage: globals_pkg